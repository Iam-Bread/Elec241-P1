-- A library clause declares a name as a library.  It 
-- does not create the library; it simply forward declares 
-- it. 
LIBRARY ieee;
USE ieee.std_logic_1164.all;
--USE ieee.std_logic_arith.all;
USE ieee.numeric_std.all;

entity SERVO is
	generic
	(
        -- Constants
		DATA_WIDTH	: integer  := 12;
		MAX_ANGLE	: integer  := 3018
	);
	port
	(
		-- Inputs
		STATE : in std_logic; --1 is on, 0 is off
		SETANGLE : in  std_logic_vector(DATA_WIDTH-1 DOWNTO 0);

		--optical encoder inputs
		OPTOA : in std_logic;	
		OPTOB : in std_logic;

        reset : in  std_logic;

		-- Outputs
		--outputs connected to hbridge to control motor
		MOTORA : out std_logic;
		MOTORB : out std_logic;

		ANGLE : out std_logic_vector(DATA_WIDTH DOWNTO 0)
	);
end SERVO;

architecture logic of SERVO is
	signal countA : std_logic_vector(DATA_WIDTH DOWNTO 0) :=(others => '0');
	signal countB : std_logic_vector(DATA_WIDTH DOWNTO 0) :=(others => '0');
	signal count : std_logic_vector(DATA_WIDTH DOWNTO 0) :=(others => '0');

begin
	ANGLE <= count;
	count<= std_logic_vector(unsigned(countA) + unsigned(countB));
	process(STATE,clk,reset)    --sensitivity list
	begin
		if(reset = '0')then		--asynchronous reset to default values
			--count <= (others=>'0') ;
			MOTORA <= '0';
			MOTORB <= '0';
		elsif(STATE = '1')then
			if(to_integer(unsigned(SETANGLE)) <= MAX_ANGLE)then	--check if angle is valid
				if(count = SETANGLE)then
					MOTORA <= '0';
					MOTORB <= '0';
				elsif(unsigned(SETANGLE) > unsigned(count))then	--check what direction to go 
					MOTORA <= '1';			--go Clockwise
					MOTORB <= '0';
				elsif(unsigned(SETANGLE) < unsigned(count))then
					MOTORA <= '0';			--go anticlockwise
					MOTORB <= '1';
				end if;
			end if;
		end if;
	end process;

	counterA: process(OPTOA)	
	begin	
		--there are 3 pulses for every 1 revolution of the motor shaft
		--as the gearbox is 1006:1 there is 3018 pulses per revolution of the output shaft

		if(rising_edge(OPTOA))then	--wait for rising edge of A
			if(unsigned(SETANGLE) > unsigned(count))then
				countA <= std_logic_vector(unsigned(countA) + 1);		--increment the count value
			else 
				countA <= std_logic_vector(unsigned(countA) - 1);		--decrement the count value
			end if;
		end if;

	end process counterA;

	counterB: process(OPTOB)	
	begin	
		--there are 3 pulses for every 1 revolution of the motor shaft
		--as the gearbox is 1006:1 there is 3018 pulses per revolution of the output shaft
		if(rising_edge(OPTOB))then
				if(unsigned(SETANGLE) > unsigned(count))then
					countB <= std_logic_vector(unsigned(countB) + 1);		--increment the count value
				else 
					countB <= std_logic_vector(unsigned(countB) - 1);		--decrement the count value
				end if;
		end if;	
	end process counterB;
end logic;